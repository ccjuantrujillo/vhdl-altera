library verilog;
use verilog.vl_types.all;
entity Multiplexor4_vlg_vec_tst is
end Multiplexor4_vlg_vec_tst;
