library verilog;
use verilog.vl_types.all;
entity Multiplexor_vlg_vec_tst is
end Multiplexor_vlg_vec_tst;
