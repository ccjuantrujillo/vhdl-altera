library verilog;
use verilog.vl_types.all;
entity compuertaAND_vlg_vec_tst is
end compuertaAND_vlg_vec_tst;
