library verilog;
use verilog.vl_types.all;
entity Altera3_vlg_vec_tst is
end Altera3_vlg_vec_tst;
