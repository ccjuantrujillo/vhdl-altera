library verilog;
use verilog.vl_types.all;
entity Alu2_vlg_vec_tst is
end Alu2_vlg_vec_tst;
