library verilog;
use verilog.vl_types.all;
entity Sumador4Bits_vlg_vec_tst is
end Sumador4Bits_vlg_vec_tst;
