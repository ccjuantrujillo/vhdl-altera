library verilog;
use verilog.vl_types.all;
entity MedioSumador_vlg_vec_tst is
end MedioSumador_vlg_vec_tst;
