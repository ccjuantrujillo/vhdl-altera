library verilog;
use verilog.vl_types.all;
entity Tutorial2_vlg_vec_tst is
end Tutorial2_vlg_vec_tst;
