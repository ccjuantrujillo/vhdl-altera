
module cpu (
	clk_clk);	

	input		clk_clk;
endmodule
