library verilog;
use verilog.vl_types.all;
entity Decoder3_6_vlg_vec_tst is
end Decoder3_6_vlg_vec_tst;
