library verilog;
use verilog.vl_types.all;
entity MedioSumador_vlg_check_tst is
    port(
        cout            : in     vl_logic;
        f               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end MedioSumador_vlg_check_tst;
